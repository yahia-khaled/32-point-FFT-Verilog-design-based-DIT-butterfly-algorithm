module Twiddle_factor_imag_ROM #(parameter WIDTH = 16)(
	input 	wire 			[2:0]				address,
	output	wire	signed	[WIDTH*16-1:0]		Twiddle_factors
);

reg			[255:0]			Twiddle_factor_ROM;


always @(*) begin
	Twiddle_factor_ROM = 0;
		case (address)
			3'b000: Twiddle_factor_ROM = 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			3'b001:	Twiddle_factor_ROM = 256'b1111111100000000000000000000000011111111000000000000000000000000111111110000000000000000000000001111111100000000000000000000000011111111000000000000000000000000111111110000000000000000000000001111111100000000000000000000000011111111000000000000000000000000;
			3'b010:	Twiddle_factor_ROM = 256'b1111111101001011111111110000000011111111010010110000000000000000111111110100101111111111000000001111111101001011000000000000000011111111010010111111111100000000111111110100101100000000000000001111111101001011111111110000000011111111010010110000000000000000;
			3'b011:	Twiddle_factor_ROM = 256'b1111111110011110111111110100101111111111000100111111111100000000111111110001001111111111010010111111111110011110000000000000000011111111100111101111111101001011111111110001001111111111000000001111111100010011111111110100101111111111100111100000000000000000;
			3'b100:	Twiddle_factor_ROM = 256'b1111111111001110111111111001111011111111011100101111111101001011111111110010101111111111000100111111111100000101111111110000000011111111000001011111111100010011111111110010101111111111010010111111111101110010111111111001111011111111110011100000000000000000;
			default : Twiddle_factor_ROM = 0;
		endcase
end

assign Twiddle_factors = Twiddle_factor_ROM;

endmodule