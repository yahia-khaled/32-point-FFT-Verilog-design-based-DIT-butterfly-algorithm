module Twiddle_factor_real_ROM #(parameter WIDTH = 16)(
	input 	wire 				[2:0]		address,
	output	wire	signed		[WIDTH*16-1:0]		Twiddle_factors
);


reg			[255:0]			Twiddle_factor_ROM;

always @(*) begin
	Twiddle_factor_ROM = 0;
		case (address)
			3'b000: Twiddle_factor_ROM = 256'b0000000100000000000000010000000000000001000000000000000100000000000000010000000000000001000000000000000100000000000000010000000000000001000000000000000100000000000000010000000000000001000000000000000100000000000000010000000000000001000000000000000100000000;
			3'b001:	Twiddle_factor_ROM = 256'b0000000000000000000000010000000000000000000000000000000100000000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000100000000;
			3'b010:	Twiddle_factor_ROM = 256'b1111111101001011000000000000000000000000101101010000000100000000111111110100101100000000000000000000000010110101000000010000000011111111010010110000000000000000000000001011010100000001000000001111111101001011000000000000000000000000101101010000000100000000;
			3'b011:	Twiddle_factor_ROM = 256'b1111111100010011111111110100101111111111100111100000000000000000000000000110001000000000101101010000000011101101000000010000000011111111000100111111111101001011111111111001111000000000000000000000000001100010000000001011010100000000111011010000000100000000;
			3'b100:	Twiddle_factor_ROM = 256'b1111111100000101111111110001001111111111001010111111111101001011111111110111001011111111100111101111111111001110000000000000000000000000001100100000000001100010000000001000111000000000101101010000000011010101000000001110110100000000111110110000000100000000;
			default : Twiddle_factor_ROM = 0;
		endcase
end

assign Twiddle_factors = Twiddle_factor_ROM;

endmodule